package delay_pkg is
    type array_8 is array (7 downto 0) of std_logic_vector(7 downto 0);
end package delay_pkg;

